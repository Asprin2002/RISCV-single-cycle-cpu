//CPU模块
module CPU(
	input wire clk,
	input wire rst,

	output wire [31:0] cur_pc_for_simulator,
	output wire [31:0] regfile_for_simulator[31:0]
);



endmodule